library verilog;
use verilog.vl_types.all;
entity core_tb_v_unit is
end core_tb_v_unit;
