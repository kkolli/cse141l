library verilog;
use verilog.vl_types.all;
entity data_mem_v_unit is
end data_mem_v_unit;
