library verilog;
use verilog.vl_types.all;
entity core_v_unit is
end core_v_unit;
