library verilog;
use verilog.vl_types.all;
entity definitions_v_unit is
end definitions_v_unit;
