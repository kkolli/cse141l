library verilog;
use verilog.vl_types.all;
entity alu_v_unit is
end alu_v_unit;
