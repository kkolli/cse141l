library verilog;
use verilog.vl_types.all;
entity instr_mem_v_unit is
end instr_mem_v_unit;
