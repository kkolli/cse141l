library verilog;
use verilog.vl_types.all;
entity cl_decode_v_unit is
end cl_decode_v_unit;
